module clock_div3(input clock_in,
			       input reset_n,
			       output clock_out);
	
	// Internal variables for the FFs
	reg qa, qb, qc;

	// Flip-flops A/B - positive clock edge
	always @(posedge clock_in or negedge reset_n)
	begin
	    if(!reset_n) begin
		    qa <= 1'b0;
			qb <= 1'b0;
	    end else begin
            qa <= (~qa) & (~qb);
            qb <= qa;
        end
	end
	
	// Flip-flop C - negative clock edge
	always @(negedge clock_in or negedge reset_n)
	begin
	    if(!reset_n)
		    qc <= 1'b0;
	    else
            qc <= qb;	
	end

    // Make the final OR gate (makes 50% duty cycle)
	assign clock_out = qb | qc;

endmodule