module hello_world();

	initial begin
	$display("\n\t My name is Imad and I start the course today! \n");
	end
endmodule